module testbench();
  input wire;
